package apb_master_package;
import uvm_pkg::*;
`include "uvm_macros.svh"
`include "apb_master_config.sv"
`include "apb_master_transaction.sv"
`include "apb_master_sequence.sv"
`include "apb_master_driver.sv"
`include "apb_master_monitor.sv"
`include "apb_master_sequencer.sv"
`include "apb_master_agent.sv"
`include "apb_master_scoreboard.sv"
`include "apb_master_environment.sv"
`include "apb_master_test.sv"
endpackage

