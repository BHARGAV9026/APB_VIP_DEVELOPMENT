`define ADDR_WIDTH 32
`define DATA_WIDTH 32
`define MEM_DEPTH 255
`define MAX_WAIT 5
