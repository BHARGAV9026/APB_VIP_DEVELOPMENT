`define DATA_WIDTH 32
`define ADDR_WIDTH 32
`define VALID_ADDR 255
